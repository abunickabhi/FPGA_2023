--import std_logic from the IEEE library
library ieee;
use ieee.std_logic_1164.all;

--ENTITY DECLARATION: name, inputs, outputs
entity not_button is
   port( inPort  : in std_logic;
         outPort : out std_logic);
end not_button;

--FUNCTIONAL DESCRIPTION: how the Inverter works
architecture func of not_button is
begin
   outPort <= not inPort;
end func;